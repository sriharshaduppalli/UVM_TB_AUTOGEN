interface simple_dut_if;
// input  clk
  logic  clk;
// input  rst_n
  logic  rst_n;
// input [7:0] in_data
  logic [[7:0]]  in_data;
// output  reg
  logic  reg;
// output  valid
  logic  valid;
endinterface